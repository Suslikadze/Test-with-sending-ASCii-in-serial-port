library ieee;

use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

Entity Serial is
Port(
    clk         : IN std_logic;
    